library verilog;
use verilog.vl_types.all;
entity tateti_vlg_check_tst is
    port(
        cont            : in     vl_logic;
        z               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end tateti_vlg_check_tst;
