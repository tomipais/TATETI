library verilog;
use verilog.vl_types.all;
entity bloqueador_vlg_vec_tst is
end bloqueador_vlg_vec_tst;
