library verilog;
use verilog.vl_types.all;
entity contador2000_vlg_vec_tst is
end contador2000_vlg_vec_tst;
