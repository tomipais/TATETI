library verilog;
use verilog.vl_types.all;
entity antirebote_vlg_vec_tst is
end antirebote_vlg_vec_tst;
