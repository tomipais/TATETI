library verilog;
use verilog.vl_types.all;
entity salidaserie_vlg_check_tst is
    port(
        sr_out          : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end salidaserie_vlg_check_tst;
