library verilog;
use verilog.vl_types.all;
entity contador_384_vlg_vec_tst is
end contador_384_vlg_vec_tst;
