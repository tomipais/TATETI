library verilog;
use verilog.vl_types.all;
entity infoleds_vlg_check_tst is
    port(
        senal           : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end infoleds_vlg_check_tst;
