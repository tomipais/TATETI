-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Mon Dec 01 17:49:15 2025

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY maqpulso IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        x : IN STD_LOGIC := '0';
        L : OUT STD_LOGIC
    );
END maqpulso;

ARCHITECTURE BEHAVIOR OF maqpulso IS
    TYPE type_fstate IS (uno,cero,ceroeterno);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,x)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= cero;
            L <= '0';
        ELSE
            L <= '0';
            CASE fstate IS
                WHEN uno =>
                    IF ((x = '1')) THEN
                        reg_fstate <= ceroeterno;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= uno;
                    END IF;

                    L <= '1';
                WHEN cero =>
                    IF ((x = '1')) THEN
                        reg_fstate <= uno;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= cero;
                    END IF;

                    L <= '0';
                WHEN ceroeterno =>
                    IF ((x = '1')) THEN
                        reg_fstate <= ceroeterno;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= ceroeterno;
                    END IF;

                    L <= '0';
                WHEN OTHERS => 
                    L <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
