library verilog;
use verilog.vl_types.all;
entity muxgrande_vlg_vec_tst is
end muxgrande_vlg_vec_tst;
