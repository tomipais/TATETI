library verilog;
use verilog.vl_types.all;
entity salidaserie_vlg_sample_tst is
    port(
        clk             : in     vl_logic;
        data_in         : in     vl_logic_vector(383 downto 0);
        enable          : in     vl_logic;
        load            : in     vl_logic;
        reset           : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end salidaserie_vlg_sample_tst;
