library verilog;
use verilog.vl_types.all;
entity infoleds_vlg_vec_tst is
end infoleds_vlg_vec_tst;
