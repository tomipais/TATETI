library verilog;
use verilog.vl_types.all;
entity botonera_vlg_vec_tst is
end botonera_vlg_vec_tst;
