library verilog;
use verilog.vl_types.all;
entity salidaserie_vlg_vec_tst is
end salidaserie_vlg_vec_tst;
