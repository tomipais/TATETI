library verilog;
use verilog.vl_types.all;
entity tateti_vlg_vec_tst is
end tateti_vlg_vec_tst;
