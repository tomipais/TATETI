-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Thu Nov 13 17:33:45 2025

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY tateti IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        x : IN STD_LOGIC := '0';
        T : IN STD_LOGIC := '0';
        z : OUT STD_LOGIC;
        cont : OUT STD_LOGIC
    );
END tateti;

ARCHITECTURE BEHAVIOR OF tateti IS
    TYPE type_fstate IS (ceroestable,unoestable,preguntauno,preguntacero);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
    SIGNAL reg_z : STD_LOGIC := '0';
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,x,T,reg_z)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= unoestable;
            reg_z <= '0';
            z <= '0';
            cont <= '0';
        ELSE
            reg_z <= '0';
            cont <= '0';
            z <= '0';
            CASE fstate IS
                WHEN ceroestable =>
                    IF ((x = '0')) THEN
                        reg_fstate <= ceroestable;
                    ELSIF ((x = '1')) THEN
                        reg_fstate <= preguntacero;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= ceroestable;
                    END IF;

                    cont <= '0';

                    reg_z <= '0';
                WHEN unoestable =>
                    IF ((x = '1')) THEN
                        reg_fstate <= unoestable;
                    ELSIF ((x = '0')) THEN
                        reg_fstate <= preguntauno;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= unoestable;
                    END IF;

                    cont <= '0';

                    reg_z <= '1';
                WHEN preguntauno =>
                    IF ((T = '0')) THEN
                        reg_fstate <= preguntauno;
                    ELSIF (((T = '1') AND (x = '0'))) THEN
                        reg_fstate <= ceroestable;
                    ELSIF (((T = '1') AND (x = '1'))) THEN
                        reg_fstate <= unoestable;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= preguntauno;
                    END IF;

                    cont <= '1';

                    reg_z <= '1';
                WHEN preguntacero =>
                    IF ((T = '0')) THEN
                        reg_fstate <= preguntacero;
                    ELSIF (((T = '1') AND (x = '0'))) THEN
                        reg_fstate <= ceroestable;
                    ELSIF (((T = '1') AND (x = '1'))) THEN
                        reg_fstate <= unoestable;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= preguntacero;
                    END IF;

                    cont <= '1';

                    reg_z <= '0';
                WHEN OTHERS => 
                    reg_z <= 'X';
                    cont <= 'X';
                    report "Reach undefined state";
            END CASE;
            z <= reg_z;
        END IF;
    END PROCESS;
END BEHAVIOR;
