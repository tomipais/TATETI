-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Mon Nov 10 16:29:32 2025

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY botonera IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        x0 : IN STD_LOGIC := '0';
        x1 : IN STD_LOGIC := '0';
        x2 : IN STD_LOGIC := '0';
        x3 : IN STD_LOGIC := '0';
        Z0 : out std_logic;
		  Z1 : out std_logic;
		  Z2 : out std_logic;
		  Z3 : out std_logic	  
    );
END botonera;

ARCHITECTURE BEHAVIOR OF botonera IS
    TYPE type_fstate IS (In2,In0,In3,In1,fijo0,fijo1,fijo2,fijo3);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
	 signal Z : STD_LOGIC_VECTOR(0 TO 3);
BEGIN
    PROCESS (clock,reset,reg_fstate)
    BEGIN
        IF (reset='1') THEN
            fstate <= In0;
        ELSIF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,x0,x1,x2,x3)
    BEGIN
        Z <= "0000";
        CASE fstate IS
            WHEN In2 =>
                IF (((((x0 = '0') AND (x1 = '0')) AND (x2 = '1')) AND (x3 = '0'))) THEN
                    reg_fstate <= fijo2;
                ELSIF ((NOT(x2) = '1')) THEN
                    reg_fstate <= In3;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= In2;
                END IF;

                Z <= "0100";
            WHEN In0 =>
                IF (((((x0 = '1') AND (x1 = '0')) AND (x2 = '0')) AND (x3 = '0'))) THEN
                    reg_fstate <= fijo0;
                ELSIF ((NOT(x0) = '1')) THEN
                    reg_fstate <= In1;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= In0;
                END IF;

                Z <= "0001";
            WHEN In3 =>
                IF (((((x0 = '0') AND (x1 = '0')) AND (x2 = '0')) AND (x3 = '1'))) THEN
                    reg_fstate <= fijo3;
                ELSIF ((NOT(x3) = '1')) THEN
                    reg_fstate <= In0;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= In3;
                END IF;

                Z <= "1000";
            WHEN In1 =>
                IF (((((x0 = '0') AND (x1 = '1')) AND (x2 = '0')) AND (x3 = '0'))) THEN
                    reg_fstate <= fijo1;
                ELSIF ((NOT(x1) = '1')) THEN
                    reg_fstate <= In2;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= In1;
                END IF;

                Z <= "0010";
            WHEN fijo0 =>
                reg_fstate <= fijo0;

                Z <= "0001";
            WHEN fijo1 =>
                reg_fstate <= fijo1;

                Z <= "0010";
            WHEN fijo2 =>
                reg_fstate <= fijo2;

                Z <= "0100";
            WHEN fijo3 =>
                reg_fstate <= fijo3;

                Z <= "1000";
            WHEN OTHERS => 
                Z <= "XXXX";
                report "Reach undefined state";
        END CASE;
    END PROCESS;
	 Z0<=Z(0);
	 Z1<=Z(1);
	 Z2<=Z(2);
	 Z3<=Z(3);
	 
END BEHAVIOR;
