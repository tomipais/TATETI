-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Mon Nov 24 22:52:11 2025

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY infoleds IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        c0 : IN STD_LOGIC := '0';
        c1 : IN STD_LOGIC := '0';
        senal : OUT STD_LOGIC
    );
END infoleds;

ARCHITECTURE BEHAVIOR OF infoleds IS
    TYPE type_fstate IS (Sig0,Sig1);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,c0,c1)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= Sig0;
            senal <= '0';
        ELSE
            senal <= '0';
            CASE fstate IS
                WHEN Sig0 =>
                    IF (((c1 = '1') AND (c0 /= '1'))) THEN
                        reg_fstate <= Sig1;
                    ELSIF (((c0 = '1') AND (c1 /= '1'))) THEN
                        reg_fstate <= Sig0;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Sig0;
                    END IF;

                    senal <= '0';
                WHEN Sig1 =>
                    IF (((c0 = '1') AND (c1 /= '1'))) THEN
                        reg_fstate <= Sig0;
                    ELSIF (((c1 = '1') AND (c0 /= '1'))) THEN
                        reg_fstate <= Sig1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Sig1;
                    END IF;

                    senal <= '1';
                WHEN OTHERS => 
                    senal <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
