-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Thu Nov 27 12:38:19 2025

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY bloqueador IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        c0 : IN STD_LOGIC := '0';
        c1 : IN STD_LOGIC := '0';
        c2 : IN STD_LOGIC := '0';
        c3 : IN STD_LOGIC := '0';
        sal0 : OUT STD_LOGIC;
        sa1 : OUT STD_LOGIC;
        sal2 : OUT STD_LOGIC;
        sal3 : OUT STD_LOGIC
    );
END bloqueador;

ARCHITECTURE BEHAVIOR OF bloqueador IS
    TYPE type_fstate IS (uno,dos,tres,block0,block1,block2,block3,cero);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reset,reg_fstate)
    BEGIN
        IF (reset='1') THEN
            fstate <= cero;
        ELSIF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,c0,c1,c2,c3)
    BEGIN
        sal0 <= '0';
        sa1 <= '0';
        sal2 <= '0';
        sal3 <= '0';
        CASE fstate IS
            WHEN uno =>
                IF (((((c0 = '0') AND (c1 = '1')) AND (c2 = '0')) AND (c3 = '0'))) THEN
                    reg_fstate <= block1;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= uno;
                END IF;

                sal2 <= '0';

                sa1 <= '1';

                sal3 <= '0';

                sal0 <= '0';
            WHEN dos =>
                IF (((((c0 = '0') AND (c1 = '0')) AND (c2 = '1')) AND (c3 = '0'))) THEN
                    reg_fstate <= block2;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= dos;
                END IF;

                sal2 <= '1';

                sa1 <= '0';

                sal3 <= '0';

                sal0 <= '0';
            WHEN tres =>
                IF (((((c0 = '1') AND (c1 = '0')) AND (c2 = '0')) AND (c3 = '1'))) THEN
                    reg_fstate <= block3;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= tres;
                END IF;

                sal2 <= '0';

                sa1 <= '0';

                sal3 <= '1';

                sal0 <= '0';
            WHEN block0 =>
                reg_fstate <= block0;

                sal0 <= '1';
            WHEN block1 =>
                reg_fstate <= block1;

                sa1 <= '1';
            WHEN block2 =>
                reg_fstate <= block2;

                sal2 <= '1';
            WHEN block3 =>
                reg_fstate <= block3;

                sal3 <= '1';
            WHEN cero =>
                IF (((((c0 = '1') AND (c1 = '0')) AND (c2 = '0')) AND (c3 = '0'))) THEN
                    reg_fstate <= block0;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= cero;
                END IF;

                sal2 <= '0';

                sa1 <= '0';

                sal3 <= '0';

                sal0 <= '1';
            WHEN OTHERS => 
                sal0 <= 'X';
                sa1 <= 'X';
                sal2 <= 'X';
                sal3 <= 'X';
                report "Reach undefined state";
        END CASE;
    END PROCESS;
END BEHAVIOR;
